
//****************************************VSCODE PLUG-IN**********************************//
//----------------------------------------------------------------------------------------
// IDE :                   VSCODE     
// VSCODE plug-in version: Verilog-Hdl-Format-2.6.20240622
// VSCODE plug-in author : Jiang Percy
//----------------------------------------------------------------------------------------
//****************************************Copyright (c)***********************************//
// Copyright(C)            Please Write Company name
// All rights reserved     
// File name:              
// Last modified Date:     2024/07/12 17:14:37
// Last Version:           V1.0
// Descriptions:           
//----------------------------------------------------------------------------------------
// Created by:             Please Write You Name 
// Created date:           2024/07/12 17:14:37
// mail      :             Please Write mail 
// Version:                V1.0
// TEXT NAME:              test2.v
// PATH:                   C:\Users\a1321\Desktop\fpga_project\cpu\user\src\test2.v
// Descriptions:           
//                         
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module test2(
    input                               clk                        ,
    input                               rst_n       ,
    output  test_out              
);
assign test_out = clk;                                  

                                                                   
                                                                   
endmodule