//****************************************VSCODE PLUG-IN**********************************//
//----------------------------------------------------------------------------------------
// IDE :                   VSCODE
// VSCODE plug-in version: Verilog-Hdl-Format-2.6.20240622
// VSCODE plug-in author : Jiang Percy
//----------------------------------------------------------------------------------------
//****************************************Copyright (c)***********************************//
// Copyright(C)            Please Write Company name
// All rights reserved
// File name:
// Last modified Date:     2024/07/14 11:19:50
// Last Version:           V1.0
// Descriptions:
//----------------------------------------------------------------------------------------
// Created by:             Please Write You Name
// Created date:           2024/07/14 11:19:50
// mail      :             Please Write mail
// Version:                V1.0
// TEXT NAME:              micro_Rom_wire.v
// PATH:                   C:\Users\a1321\Desktop\fpga_project\cpu\user\src\micro_Rom_wire.v
// Descriptions:
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module micro_Rom_wire(
        input wire [5:0]                       micro_addr,
        output wire [25:0]                   micro_op
    );
    assign micro_op = (micro_addr == 6'd0) ? 26'b00000100000000000000_000001:
                      (micro_addr == 6'd1) ? 26'b00000000000000000000_000010:
                      (micro_addr == 6'd2) ? 26'b00001000000000000100_000000:
                      (micro_addr == 6'd3) ? 26'b00000000100000100000_000000:
                      (micro_addr == 6'd4) ? 26'b00000001000000001000_000101:
                      (micro_addr == 6'd5) ? 26'b01000000000000010000_000110:
                      (micro_addr == 6'd6) ? 26'b00000000000000010000_000111:
                      (micro_addr == 6'd7) ? 26'b00000000100000010000_000000:
                      (micro_addr == 6'd8) ? 26'b00000000100101000000_000000:
                      (micro_addr == 6'd9) ? 26'b00000000001000000000_000000:
                     (micro_addr == 6'd10) ? 26'b00000000000000000010_000000:
                     (micro_addr == 6'd11) ? 26'b00010000000000100000_000000:
                     (micro_addr == 6'd12) ? 26'b00000000000000000001_000000:
                     (micro_addr == 6'd13) ? 26'b00010000000000100000_000000:
                     (micro_addr == 6'd14) ? 26'b00000000100011000000_000000:
                     (micro_addr == 6'd15) ? 26'b00000001000000001000_000000:
                     (micro_addr == 6'd16) ? 26'b10000000000000001000_010001:
                     (micro_addr == 6'd17) ? 26'b00000000000000001000_000000:
                     (micro_addr == 6'd18) ? 26'b00000000000000001000_000000:
                                             26'b00000100000000000000_000001;
endmodule
